module capture

import logger

//  TODO: document capture_region
pub fn (cap X11Capturer) capture_region(x int, y int, w int, h int) ![]u8 {
	logger.debug('capture_region start function')

	return error('not implemented yet!!!')
}
