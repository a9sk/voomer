module render

import logger

//  TODO: document init_gl_window
pub fn init_gl_window() {
	logger.debug('initializing gl window')
}

//  TODO: document draw_zoom
pub fn draw_zoom(img []u8) {
	logger.debug('draw_zoom start function')
}
