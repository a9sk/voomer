module render

import logger

pub fn init_gl_window() {
	logger.debug('initializing gl window')
}

pub fn draw_zoom(img []u8) {
	logger.debug('draw_zoom start function')
}
